module IDStage( clk , PC_i , instr );
    input clk;
    input [31:0] PC_i,instr;
    
endmodule
